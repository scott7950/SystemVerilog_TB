`ifndef __CPU_DEFINE_SV__
`define __CPU_DEFINE_SV__

typedef class cpu_transaction;
typedef mailbox #(cpu_transaction) cpu_tran_mbox;

`endif

