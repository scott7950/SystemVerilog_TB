`ifndef __PACKET_DEFINE_SV__
`define __PACKET_DEFINE_SV__

typedef class packet_transaction;
typedef mailbox #(packet_transaction) packet_tran_mbox;

`endif

